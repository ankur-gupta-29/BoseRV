module alu(
input [31:0] a,b,
input [3:0] op,
output reg [31:0] result
);
endmodule
