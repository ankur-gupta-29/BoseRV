module regfile(
input clk;
input we;
input [4:0] rs1,rs2,rd;
input [31:0] wdata;
output [31:0] rdata1,rdata2;
);
endmodule

