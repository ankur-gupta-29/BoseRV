module decode(
input [31:0] instr,
output [6:0] opcode,
output [4:0] rd,
output [2:0] funct3,
output [4:0] rs1,
output [4:0] rs2,
output [6:0] funct7,
output [31:0] imm
);


endmodule