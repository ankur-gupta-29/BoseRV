module dmem(
input clk,
input we,
input [31:0] addr,wd,
output [31:0] rd
);
endmodule;

